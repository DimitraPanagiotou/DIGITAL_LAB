`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:32:25 10/21/2020 
// Design Name: 
// Module Name:    FourDigitLEDdriver 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module FourDigitLEDdriver(rst, clk, button, an3, an2, an1, an0,
a, b, c, d, e, f, g, dp);

input clk, rst, button;
output an3, an2, an1, an0;
output a, b, c, d, e, f, g, dp;


wire new_rst,clean_btn;
wire[3:0] char;
wire[6:0] LED;

//module which synchronizes clock with reset 
//we only have posedge reset on a posedge clock
resetSynchronizer synchronizer(
		.clk(clk), 
		.rst(rst), 
		.new_rst(new_rst)
	);

//module which clean the pulse coming from the button
debouncer Debouncer(
		.rst(new_rst),
		.clk(clk),
		.noise(button),
		.clean(clean_btn)
	);
	
//module which defines the state according to a counter	
FSM mainControler(
		.clk(clk), 
		.rst(new_rst),
		.btn(clean_btn),
		.an3(an3), 
		.an2(an2), 
		.an1(an1), 
		.an0(an0), 
		.char(char)
	);	


//a simple decoder which drives the LED signals for the different char values 
LEDdecoder decoder(
		.char(char),
		.LED(LED)
	);


assign a  = LED[6];
assign b  = LED[5];
assign c  = LED[4];
assign d  = LED[3];
assign e  = LED[2];
assign f  = LED[1];
assign g  = LED[0];
assign dp = 1'b1;

endmodule
