`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:10:42 12/07/2020 
// Design Name: 
// Module Name:    bram 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module bram(clk, reset, en, address, red, green, blue);
input clk,reset,en;
input [13:0] address;
output red , green , blue;




//blockRam for red color
  RAMB16_S1 #(
      
      .INIT(1'b1),  // Value of output RAM registers at startup
      .SRVAL(1'b1), // Output value upon SSR assertion
      .WRITE_MODE("READ_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
      
		//red area
		
		.INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF), //   [0-255] binary [00000000000000 - 00000011111111]
      .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF), // [256-511] binary [00000100000000 - 00000111111111]
      .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF), // [512-767] binary [00001000000000 - 00001011111111]
      
		.INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF), //[768-1023] binary [00001100000000 - 00001111111111]
      .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[1024-1279] binary [00010000000000 - 00010011111111]
      .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[1280-1535] binary [00010100000000 - 00010111111111]
      
		.INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[1536-1791] binary [00011000000000 - 00011011111111]
      .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[1792-2047] binary [00011100000000 - 00011111111111]
      .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[2048-2303] binary [00100000000000 - 00100011111111]
      
		.INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[2304-2559] binary [00100100000000 - 00100111111111]
      .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[2560-2815] binary [00101000000000 - 00101011111111]
      .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[2816-3071] binary [00101100000000 - 00101111111111]
      
		
		//blue area
		.INIT_0C(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[3072-3327] binary [00110000000000 - 00110011111111]
      .INIT_0D(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[3328-3583] binary [00110100000000 - 00110111111111]
      .INIT_0E(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[3584-3839] binary [00111000000000 - 00111011111111]
      
		.INIT_0F(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[3840-4095] binary [00111100000000 - 00111111111111]
      .INIT_10(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[4096-4351] binary [01000000000000 - 01000011111111]
      .INIT_11(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[4352-4607] binary [01000100000000 - 01000111111111]
      
		.INIT_12(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[4608-4863] binary [01001000000000 - 01001011111111]
      .INIT_13(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[4864-5119] binary [01001100000000 - 01001111111111]
      .INIT_14(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[5120-5375] binary [01010000000000 - 01010011111111]
      
		.INIT_15(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[5376-5631] binary [01010100000000 - 01010111111111]
      .INIT_16(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[5632-5887] binary [01011000000000 - 01011011111111]
      .INIT_17(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[5888-6143] binary [01011100000000 - 01011111111111]
      
		
		//green area
		.INIT_18(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[6144-6399] binary [01100000000000 - 01100011111111]
      .INIT_19(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[6400-6655] binary [01100100000000 - 01100111111111]
      .INIT_1A(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[6656-6911] binary [01101000000000 - 01101011111111]
      
		.INIT_1B(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[6912-7167] binary [01101100000000 - 01101111111111]
      .INIT_1C(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[7168-7423] binary [01110000000000 - 01110011111111]
      .INIT_1D(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[7424-7679] binary [01110100000000 - 01110111111111]
      
		.INIT_1E(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[7680-7935] binary [01111000000000 - 01111011111111]
      .INIT_1F(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[7936-8191] binary [01111100000000 - 01111111111111]
		.INIT_20(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[8192-8447] binary [10000000000000 - 10000011111111]
      
		.INIT_21(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[8448-8703] binary [10000100000000 - 10000111111111]
      .INIT_22(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[8704-8959] binary [10001000000000 - 10001011111111]
      .INIT_23(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[8960-9215] binary [10001100000000 - 10001111111111]
      
		
		//vertical multicolor area
		//purple white light_blue black yellow
		.INIT_24(256'h0000000000003FFFFFFFFFFFFFFFFFFF_0000000000003FFFFFFFFFFFFFFFFFFF),//[9216-9471] binary [10010000000000 - 10010011111111]
      .INIT_25(256'h0000000000003FFFFFFFFFFFFFFFFFFF_0000000000003FFFFFFFFFFFFFFFFFFF),//[9472-9727] binary [10010100000000 - 10010111111111]
      .INIT_26(256'h0000000000003FFFFFFFFFFFFFFFFFFF_0000000000003FFFFFFFFFFFFFFFFFFF),//[9728-9983] binary [10011000000000 - 10011011111111]
      
		.INIT_27(256'h0000000000003FFFFFFFFFFFFFFFFFFF_0000000000003FFFFFFFFFFFFFFFFFFF),  //[9984-10239] binary [10011100000000 - 10011111111111]
      .INIT_28(256'h0000000000003FFFFFFFFFFFFFFFFFFF_0000000000003FFFFFFFFFFFFFFFFFFF), //[10240-10495] binary [10100000000000 - 10100011111111]
      .INIT_29(256'h0000000000003FFFFFFFFFFFFFFFFFFF_0000000000003FFFFFFFFFFFFFFFFFFF), //[10496-10751] binary [10100100000000 - 10100111111111]
      
		.INIT_2A(256'h0000000000003FFFFFFFFFFFFFFFFFFF_0000000000003FFFFFFFFFFFFFFFFFFF), //[10752-11007] binary [10101000000000 - 10101011111111]
      .INIT_2B(256'h0000000000003FFFFFFFFFFFFFFFFFFF_0000000000003FFFFFFFFFFFFFFFFFFF), //[11008-11263] binary [10101100000000 - 10101111111111]
      .INIT_2C(256'h0000000000003FFFFFFFFFFFFFFFFFFF_0000000000003FFFFFFFFFFFFFFFFFFF), //[11264-11519] binary [10110000000000 - 10110011111111]
      
		.INIT_2D(256'h0000000000003FFFFFFFFFFFFFFFFFFF_0000000000003FFFFFFFFFFFFFFFFFFF), //[11520-11775] binary [10110100000000 - 10110111111111]
      .INIT_2E(256'h0000000000003FFFFFFFFFFFFFFFFFFF_0000000000003FFFFFFFFFFFFFFFFFFF), //[11776-12031] binary [10111000000000 - 10111011111111]
      .INIT_2F(256'h0000000000003FFFFFFFFFFFFFFFFFFF_0000000000003FFFFFFFFFFFFFFFFFFF), //[12032-12287] binary [10111100000000 - 10111111111111]
      
		
		//memory space which is unused
		
		.INIT_30(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_31(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_32(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_33(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_34(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_35(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_36(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_37(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_38(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_39(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
      
     
   ) RED_RAMB16_S1_inst (
      .DO(red),      // 1-bit Data Output
      .ADDR(address),  // 14-bit Address Input
      .CLK(clk),    // Clock
      .DI(1'b0),      // 1-bit Data Input
      .EN(en),      // RAM Enable Input
      .SSR(reset),    // Synchronous Set/Reset Input
      .WE(1'b0)       // Write Enable Input        // Input write enable, width defined by write port depth
   );


//blockRam for green color
   RAMB16_S1 #(
      .INIT(1'b1),  // Value of output RAM registers at startup
      .SRVAL(1'b1), // Output value upon SSR assertion
      .WRITE_MODE("READ_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
      
		//red area
		
		.INIT_00(256'h00000000000000000000000000000000_00000000000000000000000000000000), //   [0-255] binary [00000000000000 - 00000011111111]
      .INIT_01(256'h00000000000000000000000000000000_00000000000000000000000000000000), // [256-511] binary [00000100000000 - 00000111111111]
      .INIT_02(256'h00000000000000000000000000000000_00000000000000000000000000000000), // [512-767] binary [00001000000000 - 00001011111111]
     
		.INIT_03(256'h00000000000000000000000000000000_00000000000000000000000000000000), //[768-1023] binary [00001100000000 - 00001111111111]
      .INIT_04(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[1024-1279] binary [00010000000000 - 00010011111111]
      .INIT_05(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[1280-1535] binary [00010100000000 - 00010111111111]
      
		.INIT_06(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[1536-1791] binary [00011000000000 - 00011011111111]
      .INIT_07(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[1792-2047] binary [00011100000000 - 00011111111111]
      .INIT_08(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[2048-2303] binary [00100000000000 - 00100011111111]
      
		.INIT_09(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[2304-2559] binary [00100100000000 - 00100111111111]
      .INIT_0A(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[2560-2815] binary [00101000000000 - 00101011111111]
      .INIT_0B(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[2816-3071] binary [00101100000000 - 00101111111111]
      
		
		//blue area
		.INIT_0C(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[3072-3327] binary [00110000000000 - 00110011111111]
      .INIT_0D(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[3328-3583] binary [00110100000000 - 00110111111111]
      .INIT_0E(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[3584-3839] binary [00111000000000 - 00111011111111]
      
		.INIT_0F(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[3840-4095] binary [00111100000000 - 00111111111111]
      .INIT_10(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[4096-4351] binary [01000000000000 - 01000011111111]
      .INIT_11(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[4352-4607] binary [01000100000000 - 01000111111111]
      
		.INIT_12(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[4608-4863] binary [01001000000000 - 01001011111111]
      .INIT_13(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[4864-5119] binary [01001100000000 - 01001111111111]
      .INIT_14(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[5120-5375] binary [01010000000000 - 01010011111111]
      
		.INIT_15(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[5376-5631] binary [01010100000000 - 01010111111111]
      .INIT_16(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[5632-5887] binary [01011000000000 - 01011011111111]
      .INIT_17(256'h00000000000000000000000000000000_00000000000000000000000000000000),//[5888-6143] binary [01011100000000 - 01011111111111]
      
		
		//green area
		.INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[6144-6399] binary [01100000000000 - 01100011111111]
      .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[6400-6655] binary [01100100000000 - 01100111111111]
      .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[6656-6911] binary [01101000000000 - 01101011111111]
      
		.INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[6912-7167] binary [01101100000000 - 01101111111111]
      .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[7168-7423] binary [01110000000000 - 01110011111111]
      .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[7424-7679] binary [01110100000000 - 01110111111111]
      
		.INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[7680-7935] binary [01111000000000 - 01111011111111]
      .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[7936-8191] binary [01111100000000 - 01111111111111]
		.INIT_20(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[8192-8447] binary [10000000000000 - 10000011111111]
      
		.INIT_21(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[8448-8703] binary [10000100000000 - 10000111111111]
      .INIT_22(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[8704-8959] binary [10001000000000 - 10001011111111]
      .INIT_23(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),//[8960-9215] binary [10001100000000 - 10001111111111]
      
		
		//MULTICOLOR area
		
		.INIT_24(256'hFFFFFFF000003FFFFFFFFFFFF0000000_FFFFFFF000003FFFFFFFFFFFF0000000),//[9216-9471] binary [10010000000000 - 10010011111111]
      .INIT_25(256'hFFFFFFF000003FFFFFFFFFFFF0000000_FFFFFFF000003FFFFFFFFFFFF0000000),//[9472-9727] binary [10010100000000 - 10010111111111]
      .INIT_26(256'hFFFFFFF000003FFFFFFFFFFFF0000000_FFFFFFF000003FFFFFFFFFFFF0000000),//[9728-9983] binary [10011000000000 - 10011011111111]
      
		.INIT_27(256'hFFFFFFF000003FFFFFFFFFFFF0000000_FFFFFFF000003FFFFFFFFFFFF0000000),  //[9984-10239] binary [10011100000000 - 10011111111111]
      .INIT_28(256'hFFFFFFF000003FFFFFFFFFFFF0000000_FFFFFFF000003FFFFFFFFFFFF0000000), //[10240-10495] binary [10100000000000 - 10100011111111]
      .INIT_29(256'hFFFFFFF000003FFFFFFFFFFFF0000000_FFFFFFF000003FFFFFFFFFFFF0000000), //[10496-10751] binary [10100100000000 - 10100111111111]
      
		.INIT_2A(256'hFFFFFFF000003FFFFFFFFFFFF0000000_FFFFFFF000003FFFFFFFFFFFF0000000), //[10752-11007] binary [10101000000000 - 10101011111111]
      .INIT_2B(256'hFFFFFFF000003FFFFFFFFFFFF0000000_FFFFFFF000003FFFFFFFFFFFF0000000), //[11008-11263] binary [10101100000000 - 10101111111111]
      .INIT_2C(256'hFFFFFFF000003FFFFFFFFFFFF0000000_FFFFFFF000003FFFFFFFFFFFF0000000), //[11264-11519] binary [10110000000000 - 10110011111111]
      
		.INIT_2D(256'hFFFFFFF000003FFFFFFFFFFFF0000000_FFFFFFF000003FFFFFFFFFFFF0000000), //[11520-11775] binary [10110100000000 - 10110111111111]
      .INIT_2E(256'hFFFFFFF000003FFFFFFFFFFFF0000000_FFFFFFF000003FFFFFFFFFFFF0000000), //[11776-12031] binary [10111000000000 - 10111011111111]
      .INIT_2F(256'hFFFFFFF000003FFFFFFFFFFFF0000000_FFFFFFF000003FFFFFFFFFFFF0000000), //[12032-12287] binary [10111100000000 - 10111111111111]
      
		
		//memory space which is unused
		
		.INIT_30(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_31(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_32(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_33(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_34(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_35(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_36(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_37(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_38(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_39(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
      
     
   ) GREEN_RAMB16_S1_inst (
      .DO(green),      // 1-bit Data Output
      .ADDR(address),  // 14-bit Address Input
      .CLK(clk),    // Clock
      .DI(1'b0),      // 1-bit Data Input
      .EN(en),      // RAM Enable Input
      .SSR(reset),    // Synchronous Set/Reset Input
      .WE(1'b0)       // Write Enable Input        // Input write enable, width defined by write port depth
   );

//blockRam for blue color
   RAMB16_S1 #(
      .INIT(1'b1),  // Value of output RAM registers at startup
      .SRVAL(1'b1), // Output value upon SSR assertion
      .WRITE_MODE("READ_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
      
		//red area
		
		.INIT_00(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_01(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_02(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      
		.INIT_03(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_04(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_05(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      
		.INIT_06(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_07(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_08(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      
		.INIT_09(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_0A(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_0B(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      
		
		//blue area
		.INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      
		.INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      
		.INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      
		.INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      
		
		//green area
		.INIT_18(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_19(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_1A(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      
		.INIT_1B(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_1C(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_1D(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      
		.INIT_1E(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_1F(256'h00000000000000000000000000000000_00000000000000000000000000000000),
		.INIT_20(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      
		.INIT_21(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_22(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      .INIT_23(256'h00000000000000000000000000000000_00000000000000000000000000000000),
      
		
		//multicolor area
		
		.INIT_24(256'hFFFFFFF0000000000003FFFFFFFFFFFF_FFFFFFF0000000000003FFFFFFFFFFFF),
      .INIT_25(256'hFFFFFFF0000000000003FFFFFFFFFFFF_FFFFFFF0000000000003FFFFFFFFFFFF),
      .INIT_26(256'hFFFFFFF0000000000003FFFFFFFFFFFF_FFFFFFF0000000000003FFFFFFFFFFFF),
      
		.INIT_27(256'hFFFFFFF0000000000003FFFFFFFFFFFF_FFFFFFF0000000000003FFFFFFFFFFFF),
      .INIT_28(256'hFFFFFFF0000000000003FFFFFFFFFFFF_FFFFFFF0000000000003FFFFFFFFFFFF),
      .INIT_29(256'hFFFFFFF0000000000003FFFFFFFFFFFF_FFFFFFF0000000000003FFFFFFFFFFFF),
      
		.INIT_2A(256'hFFFFFFF0000000000003FFFFFFFFFFFF_FFFFFFF0000000000003FFFFFFFFFFFF),
      .INIT_2B(256'hFFFFFFF0000000000003FFFFFFFFFFFF_FFFFFFF0000000000003FFFFFFFFFFFF),
      .INIT_2C(256'hFFFFFFF0000000000003FFFFFFFFFFFF_FFFFFFF0000000000003FFFFFFFFFFFF),
      
		.INIT_2D(256'hFFFFFFF0000000000003FFFFFFFFFFFF_FFFFFFF0000000000003FFFFFFFFFFFF),
      .INIT_2E(256'hFFFFFFF0000000000003FFFFFFFFFFFF_FFFFFFF0000000000003FFFFFFFFFFFF),
      .INIT_2F(256'hFFFFFFF0000000000003FFFFFFFFFFFF_FFFFFFF0000000000003FFFFFFFFFFFF),
      
		
		//memory space which is unused
		
		.INIT_30(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_31(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_32(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_33(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_34(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_35(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_36(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_37(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_38(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_39(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_3F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
     
   ) BLUE_RAMB16_S1_inst (
      .DO(blue),      // 1-bit Data Output
      .ADDR(address),  // 14-bit Address Input
      .CLK(clk),    // Clock
      .DI(1'b0),      // 1-bit Data Input
      .EN(en),      // RAM Enable Input
      .SSR(reset),    // Synchronous Set/Reset Input
      .WE(1'b0)       // Write Enable Input        // Input write enable, width defined by write port depth
   );




endmodule
